library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

entity instr_mem is
	port (
			pc: in std_logic_vector(15 downto 0);
			instruction: out  std_logic_vector(15 downto 0)
		  );
end;

architecture behav of instr_mem is
type i_mem is array (0 to 66000) of std_logic_vector(15 downto 0);
signal mem: i_mem := (others => (others => '1'));


begin


mem<=( "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000011000110000",--Add r3, r0,r6
		 "0100100110000010",--LOAD "r4",(r6)2 < stall.
		 ------------------NOP will come-------------------
		 "0000010101100010",--ADC r2,r5,"r4"
		 "0000001100100000",--Add r1, r4,r4
		 "0000010100100000",--Add r2, r4,r4
		 "0000011101110000",--Add r3, r5,r6
		 --"0000010101100010",--ADC r2,r5,"r4"
		 "0000010101110010",--ADC r2,r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000100011110000",--Add r4, "r3",r6 < forward 2nd layer.
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add "r3", r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000100101011000",--Add r4, r5,"r3" < forward 2nd layer.
		 "0000001101110000",--Add r1, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "0010001101110000",--Nnd r1, r5,r6 		
		 "0000001001000000",
		 "0000001000000000",
		 "0000001000001000",
		 
		 "0011001000000000",
		 "0000001000000000",		 
		 "0000001010011000",
		 "0000011010001000",
		 "0000011001010000",
		 "0000011001010000",
		 "0000011001010000",
		 
		 "0010100011001000",
		 "0000100010011000",
		 "0000100010011000",
		 "0000100010011000",
		 "0000100010011000",
		 "0000100010011000",
		 
		 "1100010011000000",
		 
		 "0000000000000000",
		 "0000100010011000",
		 "1001001101001010",
		 "0000110010011000",
		 "0000110010011000",
		 "0000110010011000",
		 
		 --FOR JAL
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "1000000000001001",--JAL r0, 9
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "0010001101110000",--Nnd r1, r5,r6
		 "0000001001000000",
		 "0000001000000000",
		 "0000001000001000",
		 "0011001000000000",--<-JUMP HERE
		 "0000001000000000",
		 
		 --FOR JLR
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "1001110101000000",--JLR r6, r5
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "0010001101110000",--Nnd r1, r5,r6 --<-jump here
		 "0000001001000000",
		 "0000001000000000",
		 "0000001000001000",
		 
		 --FOR BEQ
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "1100110101001101",--BEQ r6, r5, 13
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "0010001101110000",--Nnd r1, r5,r6 
		 "0000001001000000",
		 "0000001000000000",
		 "0000001000001000",
		 
		 "0011001000000000",
		 "0000001000000000",		 
		 "0000001010011000",
		 "0000011010001000",
		 "0000011001010000",--<-jump here
		 
		 -- forwarding logic 2 layer only ADD & NAND
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add "r3", r5,r6
		 "0000100011110000",--Add r4, "r3",r6 < forward.
		 "0000010101110000",--Add "r2", r5,r6
		 "0000011101010000",--Add r3, r5,"r2" < forward.
		 "0000011101110000",--Add "r3", r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000100011110000",--Add r4, "r3",r6 < forward 2nd layer.
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add "r3", r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000100101011000",--Add r4, r5,"r3" < forward 2nd layer.
		 "0000001101110000",--Add r1, r5,r6
		 "0000100101110000",--Add r4, r5,r6
		 "0010001101110000",--Nnd r1, r5,r6 
		 
		-- LOAD + stall + forwarding + ADC {image saved}
		-- (carry is passes when load, no stall, 
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011000110000",--Add r3, r0,r6
		 "0100100110000010",--LOAD "r4",(r6)2 < stall.
		 "0000010101100010",--ADC r2,r5,"r4"
		 "0000001101110000",--Add r1, r5,r6
		 "0000010101110000",--Add r2, r5,r6
		 "0000011101110000",--Add r3, r5,r6
		
		
		 "0000110010011000",
		 "0000110010011000",
		 "0000110010011000",
		 "0000110010011111",
		 "0000110010011000",
		 "0000110010011000",
		 "0000110010011000",
		 "0000110010011000",
		 "0000110010011000",
		 "0000110010011000",
		 others => (others => '1')
		);
instruction <= mem(to_integer(unsigned(pc)));

end behav;